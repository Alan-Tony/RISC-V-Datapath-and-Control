library verilog;
use verilog.vl_types.all;
entity WB_TB is
end WB_TB;
