library verilog;
use verilog.vl_types.all;
entity ALU_TopLevel_TB is
end ALU_TopLevel_TB;
