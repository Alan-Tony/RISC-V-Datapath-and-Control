library verilog;
use verilog.vl_types.all;
entity ALU_1b_Ordinary_TB is
end ALU_1b_Ordinary_TB;
