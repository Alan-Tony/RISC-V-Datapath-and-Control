library verilog;
use verilog.vl_types.all;
entity fullAdder_TB is
end fullAdder_TB;
