library verilog;
use verilog.vl_types.all;
entity ID_and_RF_TB is
end ID_and_RF_TB;
