library verilog;
use verilog.vl_types.all;
entity Memory_TB is
end Memory_TB;
