
module MyInverter (A, B);
  
  input A;
  output B;
  
  not M1(B, A);

endmodule
