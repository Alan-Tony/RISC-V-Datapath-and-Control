library verilog;
use verilog.vl_types.all;
entity Data_Memory_TB is
end Data_Memory_TB;
