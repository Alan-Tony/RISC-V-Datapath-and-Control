library verilog;
use verilog.vl_types.all;
entity signextendtestbench is
end signextendtestbench;
