library verilog;
use verilog.vl_types.all;
entity mux4to1_TB is
end mux4to1_TB;
