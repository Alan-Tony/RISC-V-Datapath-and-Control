library verilog;
use verilog.vl_types.all;
entity exec_tb is
end exec_tb;
