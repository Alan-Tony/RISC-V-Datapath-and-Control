library verilog;
use verilog.vl_types.all;
entity Pipeline is
end Pipeline;
