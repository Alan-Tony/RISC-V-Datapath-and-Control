library verilog;
use verilog.vl_types.all;
entity IF_Testbench is
end IF_Testbench;
